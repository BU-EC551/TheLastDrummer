`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:23:13 03/23/2015 
// Design Name: 
// Module Name:    sync 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module vgasync(vga_h_sync, vga_v_sync, inDisplayArea, CounterX, CounterY,pixel_clk);
input pixel_clk;
output vga_h_sync, vga_v_sync;
output inDisplayArea;
output reg[9:0] CounterX;
output reg [8:0] CounterY;

wire CounterXmaxed = (CounterX==10'h2FF);

always @(posedge pixel_clk)
if(CounterXmaxed)
	CounterX <= 0;
else
	CounterX <= CounterX + 1'b1;

always @(posedge pixel_clk)
if(CounterXmaxed) CounterY <= CounterY + 1'b1;

reg	vga_HS, vga_VS;
always @(posedge pixel_clk)
begin
	vga_HS <= (CounterX[9:4]==6'h2D); // change this value to move the display horizontally
	vga_VS <= (CounterY==500); // change this value to move the display vertically
end

reg inDisplayArea;
always @(posedge pixel_clk)
if(inDisplayArea==0)
	inDisplayArea <= (CounterXmaxed) && (CounterY<480);
else
	inDisplayArea <= !(CounterX==639);
	
assign vga_h_sync = ~vga_HS;
assign vga_v_sync = ~vga_VS;

endmodule

