`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:11:02 04/28/2015 
// Design Name: 
// Module Name:    keydetect 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module keydetect(input [11:0]xaxis,yaxis,input TP_DCLK,output reg [3:0]key
    );

always@
endmodule
